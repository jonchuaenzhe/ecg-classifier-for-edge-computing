`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 27.01.2022 17:50:18
// Design Name: 
// Module Name: Data_RAM
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module CONV1D_3rd_RAM
    #(
        Bit_width = 16,
        RAM_Depth = 512
    )
    (
        // Input
        input CLK,
        input Enable,
        input [4:0] Depth,
        input [3:0] Width,

        // Output
        output reg signed [Bit_width - 1 : 0] data_out_0,
        output reg signed [Bit_width - 1 : 0] data_out_1,
        output reg signed [Bit_width - 1 : 0] data_out_2,
        output reg signed [Bit_width - 1 : 0] data_out_3
    );

    // RAM reg creation
    (* ROM_STYLE="BLOCK"*) reg signed [Bit_width - 1 : 0] RAM_0 [0 : RAM_Depth - 1];
    (* ROM_STYLE="BLOCK"*) reg signed [Bit_width - 1 : 0] RAM_1 [0 : RAM_Depth - 1];
    (* ROM_STYLE="BLOCK"*) reg signed [Bit_width - 1 : 0] RAM_2 [0 : RAM_Depth - 1];
    (* ROM_STYLE="BLOCK"*) reg signed [Bit_width - 1 : 0] RAM_3 [0 : RAM_Depth - 1];

    // RAM Address
    wire [8:0] ADDR = (Width << 5) + Depth;

    always @ (negedge CLK) begin
        if (Enable) begin
            data_out_0 <= RAM_0[ADDR];
            data_out_1 <= RAM_1[ADDR];
            data_out_2 <= RAM_2[ADDR];
            data_out_3 <= RAM_3[ADDR];
        end else begin
            data_out_0 <= 0;
            data_out_1 <= 0;
            data_out_2 <= 0;
            data_out_3 <= 0;
        end
    end

    // Initialise weights
    initial begin
        RAM_0[0] = -16'd6;
        RAM_1[0] = -16'd3;
        RAM_2[0] = -16'd2;
        RAM_3[0] = -16'd3;
        RAM_0[1] = -16'd1;
        RAM_1[1] = 16'd0;
        RAM_2[1] = 16'd0;
        RAM_3[1] = 16'd0;
        RAM_0[2] = -16'd3;
        RAM_1[2] = -16'd1;
        RAM_2[2] = -16'd2;
        RAM_3[2] = 16'd0;
        RAM_0[3] = -16'd2;
        RAM_1[3] = 16'd0;
        RAM_2[3] = 16'd0;
        RAM_3[3] = 16'd0;
        RAM_0[4] = -16'd6;
        RAM_1[4] = 16'd0;
        RAM_2[4] = 16'd0;
        RAM_3[4] = 16'd0;
        RAM_0[5] = -16'd1;
        RAM_1[5] = 16'd3;
        RAM_2[5] = -16'd18;
        RAM_3[5] = -16'd22;
        RAM_0[6] = 16'd1;
        RAM_1[6] = -16'd9;
        RAM_2[6] = -16'd2;
        RAM_3[6] = -16'd1;
        RAM_0[7] = -16'd3;
        RAM_1[7] = -16'd3;
        RAM_2[7] = -16'd1;
        RAM_3[7] = 16'd2;
        RAM_0[8] = -16'd10;
        RAM_1[8] = -16'd15;
        RAM_2[8] = -16'd4;
        RAM_3[8] = -16'd2;
        RAM_0[9] = 16'd8;
        RAM_1[9] = -16'd9;
        RAM_2[9] = -16'd5;
        RAM_3[9] = -16'd3;
        RAM_0[10] = -16'd9;
        RAM_1[10] = 16'd0;
        RAM_2[10] = 16'd0;
        RAM_3[10] = 16'd0;
        RAM_0[11] = 16'd1;
        RAM_1[11] = 16'd0;
        RAM_2[11] = -16'd1;
        RAM_3[11] = 16'd3;
        RAM_0[12] = -16'd16;
        RAM_1[12] = 16'd0;
        RAM_2[12] = 16'd0;
        RAM_3[12] = 16'd0;
        RAM_0[13] = -16'd19;
        RAM_1[13] = -16'd7;
        RAM_2[13] = -16'd2;
        RAM_3[13] = -16'd3;
        RAM_0[14] = -16'd10;
        RAM_1[14] = 16'd0;
        RAM_2[14] = 16'd0;
        RAM_3[14] = 16'd0;
        RAM_0[15] = -16'd4;
        RAM_1[15] = 16'd0;
        RAM_2[15] = 16'd0;
        RAM_3[15] = 16'd0;
        RAM_0[16] = -16'd29;
        RAM_1[16] = -16'd4;
        RAM_2[16] = -16'd1;
        RAM_3[16] = 16'd1;
        RAM_0[17] = 16'd5;
        RAM_1[17] = 16'd2;
        RAM_2[17] = 16'd5;
        RAM_3[17] = -16'd4;
        RAM_0[18] = -16'd1;
        RAM_1[18] = 16'd0;
        RAM_2[18] = 16'd0;
        RAM_3[18] = 16'd1;
        RAM_0[19] = 16'd0;
        RAM_1[19] = -16'd10;
        RAM_2[19] = -16'd4;
        RAM_3[19] = -16'd4;
        RAM_0[20] = 16'd1;
        RAM_1[20] = -16'd18;
        RAM_2[20] = -16'd13;
        RAM_3[20] = 16'd1;
        RAM_0[21] = 16'd7;
        RAM_1[21] = -16'd5;
        RAM_2[21] = 16'd2;
        RAM_3[21] = -16'd1;
        RAM_0[22] = 16'd4;
        RAM_1[22] = 16'd0;
        RAM_2[22] = 16'd0;
        RAM_3[22] = 16'd0;
        RAM_0[23] = -16'd5;
        RAM_1[23] = -16'd6;
        RAM_2[23] = -16'd4;
        RAM_3[23] = -16'd4;
        RAM_0[24] = 16'd1;
        RAM_1[24] = -16'd1;
        RAM_2[24] = 16'd1;
        RAM_3[24] = 16'd2;
        RAM_0[25] = 16'd8;
        RAM_1[25] = -16'd11;
        RAM_2[25] = -16'd9;
        RAM_3[25] = -16'd4;
        RAM_0[26] = 16'd6;
        RAM_1[26] = -16'd19;
        RAM_2[26] = -16'd10;
        RAM_3[26] = -16'd1;
        RAM_0[27] = 16'd0;
        RAM_1[27] = -16'd14;
        RAM_2[27] = 16'd0;
        RAM_3[27] = 16'd2;
        RAM_0[28] = 16'd2;
        RAM_1[28] = -16'd13;
        RAM_2[28] = -16'd9;
        RAM_3[28] = 16'd0;
        RAM_0[29] = -16'd3;
        RAM_1[29] = -16'd4;
        RAM_2[29] = -16'd2;
        RAM_3[29] = -16'd2;
        RAM_0[30] = -16'd20;
        RAM_1[30] = 16'd6;
        RAM_2[30] = 16'd4;
        RAM_3[30] = -16'd2;
        RAM_0[31] = -16'd11;
        RAM_1[31] = 16'd0;
        RAM_2[31] = 16'd0;
        RAM_3[31] = 16'd0;
        RAM_0[32] = -16'd6;
        RAM_1[32] = 16'd0;
        RAM_2[32] = 16'd6;
        RAM_3[32] = -16'd27;
        RAM_0[33] = -16'd1;
        RAM_1[33] = -16'd8;
        RAM_2[33] = 16'd6;
        RAM_3[33] = -16'd30;
        RAM_0[34] = -16'd3;
        RAM_1[34] = -16'd11;
        RAM_2[34] = 16'd6;
        RAM_3[34] = -16'd31;
        RAM_0[35] = -16'd2;
        RAM_1[35] = 16'd2;
        RAM_2[35] = -16'd30;
        RAM_3[35] = 16'd3;
        RAM_0[36] = -16'd6;
        RAM_1[36] = 16'd0;
        RAM_2[36] = 16'd0;
        RAM_3[36] = 16'd0;
        RAM_0[37] = -16'd1;
        RAM_1[37] = 16'd5;
        RAM_2[37] = 16'd4;
        RAM_3[37] = 16'd8;
        RAM_0[38] = 16'd1;
        RAM_1[38] = 16'd13;
        RAM_2[38] = -16'd12;
        RAM_3[38] = -16'd7;
        RAM_0[39] = -16'd3;
        RAM_1[39] = -16'd4;
        RAM_2[39] = 16'd0;
        RAM_3[39] = -16'd39;
        RAM_0[40] = -16'd10;
        RAM_1[40] = 16'd11;
        RAM_2[40] = -16'd20;
        RAM_3[40] = 16'd6;
        RAM_0[41] = 16'd8;
        RAM_1[41] = 16'd1;
        RAM_2[41] = -16'd6;
        RAM_3[41] = -16'd23;
        RAM_0[42] = -16'd9;
        RAM_1[42] = 16'd0;
        RAM_2[42] = 16'd0;
        RAM_3[42] = 16'd0;
        RAM_0[43] = 16'd1;
        RAM_1[43] = -16'd6;
        RAM_2[43] = -16'd16;
        RAM_3[43] = -16'd24;
        RAM_0[44] = -16'd16;
        RAM_1[44] = 16'd0;
        RAM_2[44] = 16'd0;
        RAM_3[44] = 16'd0;
        RAM_0[45] = -16'd19;
        RAM_1[45] = -16'd7;
        RAM_2[45] = -16'd5;
        RAM_3[45] = -16'd18;
        RAM_0[46] = -16'd10;
        RAM_1[46] = 16'd0;
        RAM_2[46] = 16'd0;
        RAM_3[46] = 16'd0;
        RAM_0[47] = -16'd4;
        RAM_1[47] = 16'd0;
        RAM_2[47] = 16'd0;
        RAM_3[47] = 16'd0;
        RAM_0[48] = -16'd29;
        RAM_1[48] = -16'd4;
        RAM_2[48] = -16'd4;
        RAM_3[48] = 16'd3;
        RAM_0[49] = 16'd5;
        RAM_1[49] = 16'd1;
        RAM_2[49] = -16'd3;
        RAM_3[49] = -16'd22;
        RAM_0[50] = -16'd1;
        RAM_1[50] = -16'd1;
        RAM_2[50] = -16'd15;
        RAM_3[50] = -16'd34;
        RAM_0[51] = 16'd0;
        RAM_1[51] = -16'd7;
        RAM_2[51] = -16'd21;
        RAM_3[51] = 16'd3;
        RAM_0[52] = 16'd1;
        RAM_1[52] = 16'd8;
        RAM_2[52] = 16'd4;
        RAM_3[52] = 16'd1;
        RAM_0[53] = 16'd7;
        RAM_1[53] = 16'd5;
        RAM_2[53] = -16'd14;
        RAM_3[53] = -16'd16;
        RAM_0[54] = 16'd4;
        RAM_1[54] = 16'd0;
        RAM_2[54] = 16'd10;
        RAM_3[54] = -16'd30;
        RAM_0[55] = -16'd5;
        RAM_1[55] = 16'd4;
        RAM_2[55] = -16'd7;
        RAM_3[55] = -16'd10;
        RAM_0[56] = 16'd1;
        RAM_1[56] = -16'd5;
        RAM_2[56] = -16'd19;
        RAM_3[56] = -16'd14;
        RAM_0[57] = 16'd8;
        RAM_1[57] = 16'd11;
        RAM_2[57] = -16'd7;
        RAM_3[57] = -16'd22;
        RAM_0[58] = 16'd6;
        RAM_1[58] = 16'd8;
        RAM_2[58] = -16'd17;
        RAM_3[58] = -16'd18;
        RAM_0[59] = 16'd0;
        RAM_1[59] = -16'd10;
        RAM_2[59] = -16'd7;
        RAM_3[59] = 16'd1;
        RAM_0[60] = 16'd2;
        RAM_1[60] = 16'd3;
        RAM_2[60] = 16'd0;
        RAM_3[60] = -16'd9;
        RAM_0[61] = -16'd3;
        RAM_1[61] = 16'd5;
        RAM_2[61] = -16'd3;
        RAM_3[61] = -16'd8;
        RAM_0[62] = -16'd20;
        RAM_1[62] = -16'd14;
        RAM_2[62] = -16'd14;
        RAM_3[62] = -16'd20;
        RAM_0[63] = -16'd11;
        RAM_1[63] = 16'd0;
        RAM_2[63] = 16'd0;
        RAM_3[63] = 16'd0;
        RAM_0[64] = -16'd6;
        RAM_1[64] = -16'd14;
        RAM_2[64] = -16'd36;
        RAM_3[64] = -16'd18;
        RAM_0[65] = -16'd1;
        RAM_1[65] = -16'd19;
        RAM_2[65] = -16'd19;
        RAM_3[65] = -16'd5;
        RAM_0[66] = -16'd3;
        RAM_1[66] = -16'd28;
        RAM_2[66] = -16'd18;
        RAM_3[66] = 16'd8;
        RAM_0[67] = -16'd2;
        RAM_1[67] = -16'd9;
        RAM_2[67] = 16'd25;
        RAM_3[67] = -16'd15;
        RAM_0[68] = -16'd6;
        RAM_1[68] = 16'd0;
        RAM_2[68] = 16'd0;
        RAM_3[68] = 16'd0;
        RAM_0[69] = -16'd1;
        RAM_1[69] = 16'd11;
        RAM_2[69] = -16'd15;
        RAM_3[69] = -16'd25;
        RAM_0[70] = 16'd1;
        RAM_1[70] = -16'd12;
        RAM_2[70] = -16'd5;
        RAM_3[70] = -16'd9;
        RAM_0[71] = -16'd3;
        RAM_1[71] = -16'd28;
        RAM_2[71] = -16'd12;
        RAM_3[71] = -16'd4;
        RAM_0[72] = -16'd10;
        RAM_1[72] = 16'd2;
        RAM_2[72] = 16'd4;
        RAM_3[72] = 16'd7;
        RAM_0[73] = 16'd8;
        RAM_1[73] = 16'd2;
        RAM_2[73] = -16'd15;
        RAM_3[73] = -16'd8;
        RAM_0[74] = -16'd9;
        RAM_1[74] = 16'd0;
        RAM_2[74] = 16'd0;
        RAM_3[74] = 16'd0;
        RAM_0[75] = 16'd1;
        RAM_1[75] = -16'd7;
        RAM_2[75] = -16'd8;
        RAM_3[75] = -16'd14;
        RAM_0[76] = -16'd16;
        RAM_1[76] = 16'd0;
        RAM_2[76] = 16'd0;
        RAM_3[76] = 16'd0;
        RAM_0[77] = -16'd19;
        RAM_1[77] = 16'd4;
        RAM_2[77] = 16'd16;
        RAM_3[77] = 16'd5;
        RAM_0[78] = -16'd10;
        RAM_1[78] = 16'd0;
        RAM_2[78] = 16'd0;
        RAM_3[78] = 16'd0;
        RAM_0[79] = -16'd4;
        RAM_1[79] = 16'd0;
        RAM_2[79] = 16'd0;
        RAM_3[79] = 16'd0;
        RAM_0[80] = -16'd29;
        RAM_1[80] = -16'd4;
        RAM_2[80] = 16'd5;
        RAM_3[80] = 16'd20;
        RAM_0[81] = 16'd5;
        RAM_1[81] = -16'd4;
        RAM_2[81] = -16'd11;
        RAM_3[81] = -16'd6;
        RAM_0[82] = -16'd1;
        RAM_1[82] = -16'd13;
        RAM_2[82] = 16'd5;
        RAM_3[82] = -16'd5;
        RAM_0[83] = 16'd0;
        RAM_1[83] = -16'd4;
        RAM_2[83] = -16'd4;
        RAM_3[83] = 16'd5;
        RAM_0[84] = 16'd1;
        RAM_1[84] = -16'd24;
        RAM_2[84] = -16'd35;
        RAM_3[84] = 16'd18;
        RAM_0[85] = 16'd7;
        RAM_1[85] = -16'd9;
        RAM_2[85] = -16'd19;
        RAM_3[85] = -16'd6;
        RAM_0[86] = 16'd4;
        RAM_1[86] = -16'd29;
        RAM_2[86] = -16'd32;
        RAM_3[86] = -16'd7;
        RAM_0[87] = -16'd5;
        RAM_1[87] = 16'd1;
        RAM_2[87] = -16'd8;
        RAM_3[87] = -16'd1;
        RAM_0[88] = 16'd1;
        RAM_1[88] = -16'd13;
        RAM_2[88] = 16'd2;
        RAM_3[88] = -16'd16;
        RAM_0[89] = 16'd8;
        RAM_1[89] = -16'd6;
        RAM_2[89] = -16'd9;
        RAM_3[89] = -16'd12;
        RAM_0[90] = 16'd6;
        RAM_1[90] = -16'd3;
        RAM_2[90] = -16'd19;
        RAM_3[90] = 16'd1;
        RAM_0[91] = 16'd0;
        RAM_1[91] = -16'd1;
        RAM_2[91] = 16'd14;
        RAM_3[91] = -16'd5;
        RAM_0[92] = 16'd2;
        RAM_1[92] = 16'd16;
        RAM_2[92] = 16'd3;
        RAM_3[92] = -16'd2;
        RAM_0[93] = -16'd3;
        RAM_1[93] = -16'd1;
        RAM_2[93] = -16'd5;
        RAM_3[93] = -16'd19;
        RAM_0[94] = -16'd20;
        RAM_1[94] = 16'd0;
        RAM_2[94] = 16'd2;
        RAM_3[94] = 16'd5;
        RAM_0[95] = -16'd11;
        RAM_1[95] = 16'd0;
        RAM_2[95] = 16'd0;
        RAM_3[95] = 16'd0;
        RAM_0[96] = -16'd6;
        RAM_1[96] = 16'd16;
        RAM_2[96] = -16'd8;
        RAM_3[96] = -16'd9;
        RAM_0[97] = -16'd1;
        RAM_1[97] = 16'd8;
        RAM_2[97] = -16'd1;
        RAM_3[97] = 16'd7;
        RAM_0[98] = -16'd3;
        RAM_1[98] = 16'd11;
        RAM_2[98] = -16'd5;
        RAM_3[98] = 16'd12;
        RAM_0[99] = -16'd2;
        RAM_1[99] = 16'd15;
        RAM_2[99] = 16'd5;
        RAM_3[99] = 16'd1;
        RAM_0[100] = -16'd6;
        RAM_1[100] = 16'd0;
        RAM_2[100] = 16'd0;
        RAM_3[100] = 16'd0;
        RAM_0[101] = -16'd1;
        RAM_1[101] = -16'd13;
        RAM_2[101] = -16'd14;
        RAM_3[101] = -16'd26;
        RAM_0[102] = 16'd1;
        RAM_1[102] = 16'd18;
        RAM_2[102] = -16'd10;
        RAM_3[102] = -16'd21;
        RAM_0[103] = -16'd3;
        RAM_1[103] = 16'd8;
        RAM_2[103] = 16'd7;
        RAM_3[103] = 16'd7;
        RAM_0[104] = -16'd10;
        RAM_1[104] = -16'd19;
        RAM_2[104] = -16'd1;
        RAM_3[104] = -16'd9;
        RAM_0[105] = 16'd8;
        RAM_1[105] = -16'd26;
        RAM_2[105] = -16'd11;
        RAM_3[105] = 16'd2;
        RAM_0[106] = -16'd9;
        RAM_1[106] = 16'd0;
        RAM_2[106] = 16'd0;
        RAM_3[106] = 16'd0;
        RAM_0[107] = 16'd1;
        RAM_1[107] = 16'd16;
        RAM_2[107] = 16'd6;
        RAM_3[107] = -16'd3;
        RAM_0[108] = -16'd16;
        RAM_1[108] = 16'd0;
        RAM_2[108] = 16'd0;
        RAM_3[108] = 16'd0;
        RAM_0[109] = -16'd19;
        RAM_1[109] = -16'd7;
        RAM_2[109] = -16'd14;
        RAM_3[109] = 16'd6;
        RAM_0[110] = -16'd10;
        RAM_1[110] = 16'd0;
        RAM_2[110] = 16'd0;
        RAM_3[110] = 16'd0;
        RAM_0[111] = -16'd4;
        RAM_1[111] = 16'd0;
        RAM_2[111] = 16'd0;
        RAM_3[111] = 16'd0;
        RAM_0[112] = -16'd29;
        RAM_1[112] = -16'd7;
        RAM_2[112] = 16'd7;
        RAM_3[112] = -16'd11;
        RAM_0[113] = 16'd5;
        RAM_1[113] = -16'd21;
        RAM_2[113] = -16'd4;
        RAM_3[113] = -16'd4;
        RAM_0[114] = -16'd1;
        RAM_1[114] = 16'd17;
        RAM_2[114] = 16'd10;
        RAM_3[114] = 16'd11;
        RAM_0[115] = 16'd0;
        RAM_1[115] = -16'd15;
        RAM_2[115] = 16'd6;
        RAM_3[115] = -16'd4;
        RAM_0[116] = 16'd1;
        RAM_1[116] = 16'd2;
        RAM_2[116] = -16'd13;
        RAM_3[116] = -16'd7;
        RAM_0[117] = 16'd7;
        RAM_1[117] = -16'd39;
        RAM_2[117] = -16'd10;
        RAM_3[117] = 16'd9;
        RAM_0[118] = 16'd4;
        RAM_1[118] = 16'd8;
        RAM_2[118] = -16'd12;
        RAM_3[118] = -16'd1;
        RAM_0[119] = -16'd5;
        RAM_1[119] = -16'd29;
        RAM_2[119] = 16'd1;
        RAM_3[119] = -16'd3;
        RAM_0[120] = 16'd1;
        RAM_1[120] = 16'd0;
        RAM_2[120] = 16'd5;
        RAM_3[120] = -16'd1;
        RAM_0[121] = 16'd8;
        RAM_1[121] = -16'd26;
        RAM_2[121] = -16'd15;
        RAM_3[121] = -16'd1;
        RAM_0[122] = 16'd6;
        RAM_1[122] = -16'd31;
        RAM_2[122] = -16'd7;
        RAM_3[122] = -16'd4;
        RAM_0[123] = 16'd0;
        RAM_1[123] = -16'd9;
        RAM_2[123] = 16'd4;
        RAM_3[123] = 16'd6;
        RAM_0[124] = 16'd2;
        RAM_1[124] = -16'd25;
        RAM_2[124] = -16'd3;
        RAM_3[124] = 16'd1;
        RAM_0[125] = -16'd3;
        RAM_1[125] = 16'd10;
        RAM_2[125] = 16'd6;
        RAM_3[125] = -16'd24;
        RAM_0[126] = -16'd20;
        RAM_1[126] = 16'd0;
        RAM_2[126] = 16'd2;
        RAM_3[126] = -16'd18;
        RAM_0[127] = -16'd11;
        RAM_1[127] = 16'd0;
        RAM_2[127] = 16'd0;
        RAM_3[127] = 16'd0;
        RAM_0[128] = -16'd6;
        RAM_1[128] = -16'd5;
        RAM_2[128] = 16'd3;
        RAM_3[128] = -16'd1;
        RAM_0[129] = -16'd1;
        RAM_1[129] = -16'd23;
        RAM_2[129] = -16'd26;
        RAM_3[129] = 16'd8;
        RAM_0[130] = -16'd3;
        RAM_1[130] = 16'd8;
        RAM_2[130] = -16'd10;
        RAM_3[130] = 16'd25;
        RAM_0[131] = -16'd2;
        RAM_1[131] = -16'd20;
        RAM_2[131] = -16'd4;
        RAM_3[131] = -16'd27;
        RAM_0[132] = -16'd6;
        RAM_1[132] = 16'd0;
        RAM_2[132] = 16'd0;
        RAM_3[132] = 16'd0;
        RAM_0[133] = -16'd1;
        RAM_1[133] = -16'd37;
        RAM_2[133] = 16'd6;
        RAM_3[133] = 16'd0;
        RAM_0[134] = 16'd1;
        RAM_1[134] = -16'd2;
        RAM_2[134] = 16'd5;
        RAM_3[134] = -16'd1;
        RAM_0[135] = -16'd3;
        RAM_1[135] = 16'd2;
        RAM_2[135] = -16'd15;
        RAM_3[135] = 16'd20;
        RAM_0[136] = -16'd10;
        RAM_1[136] = -16'd7;
        RAM_2[136] = -16'd3;
        RAM_3[136] = -16'd2;
        RAM_0[137] = 16'd8;
        RAM_1[137] = -16'd6;
        RAM_2[137] = -16'd8;
        RAM_3[137] = 16'd5;
        RAM_0[138] = -16'd9;
        RAM_1[138] = 16'd0;
        RAM_2[138] = 16'd0;
        RAM_3[138] = 16'd0;
        RAM_0[139] = 16'd1;
        RAM_1[139] = 16'd3;
        RAM_2[139] = 16'd1;
        RAM_3[139] = -16'd13;
        RAM_0[140] = -16'd16;
        RAM_1[140] = 16'd0;
        RAM_2[140] = 16'd0;
        RAM_3[140] = 16'd0;
        RAM_0[141] = -16'd19;
        RAM_1[141] = 16'd5;
        RAM_2[141] = -16'd8;
        RAM_3[141] = -16'd16;
        RAM_0[142] = -16'd10;
        RAM_1[142] = 16'd0;
        RAM_2[142] = 16'd0;
        RAM_3[142] = 16'd0;
        RAM_0[143] = -16'd4;
        RAM_1[143] = 16'd0;
        RAM_2[143] = 16'd0;
        RAM_3[143] = 16'd0;
        RAM_0[144] = -16'd29;
        RAM_1[144] = 16'd1;
        RAM_2[144] = -16'd1;
        RAM_3[144] = 16'd0;
        RAM_0[145] = 16'd5;
        RAM_1[145] = -16'd6;
        RAM_2[145] = -16'd5;
        RAM_3[145] = 16'd2;
        RAM_0[146] = -16'd1;
        RAM_1[146] = 16'd2;
        RAM_2[146] = -16'd11;
        RAM_3[146] = -16'd8;
        RAM_0[147] = 16'd0;
        RAM_1[147] = -16'd13;
        RAM_2[147] = 16'd1;
        RAM_3[147] = -16'd6;
        RAM_0[148] = 16'd1;
        RAM_1[148] = 16'd10;
        RAM_2[148] = -16'd19;
        RAM_3[148] = 16'd14;
        RAM_0[149] = 16'd7;
        RAM_1[149] = -16'd6;
        RAM_2[149] = -16'd12;
        RAM_3[149] = 16'd14;
        RAM_0[150] = 16'd4;
        RAM_1[150] = -16'd12;
        RAM_2[150] = -16'd12;
        RAM_3[150] = 16'd4;
        RAM_0[151] = -16'd5;
        RAM_1[151] = -16'd3;
        RAM_2[151] = 16'd8;
        RAM_3[151] = 16'd15;
        RAM_0[152] = 16'd1;
        RAM_1[152] = 16'd4;
        RAM_2[152] = 16'd7;
        RAM_3[152] = -16'd18;
        RAM_0[153] = 16'd8;
        RAM_1[153] = -16'd11;
        RAM_2[153] = -16'd18;
        RAM_3[153] = 16'd10;
        RAM_0[154] = 16'd6;
        RAM_1[154] = -16'd12;
        RAM_2[154] = -16'd20;
        RAM_3[154] = 16'd18;
        RAM_0[155] = 16'd0;
        RAM_1[155] = 16'd1;
        RAM_2[155] = -16'd1;
        RAM_3[155] = 16'd5;
        RAM_0[156] = 16'd2;
        RAM_1[156] = -16'd8;
        RAM_2[156] = -16'd3;
        RAM_3[156] = -16'd8;
        RAM_0[157] = -16'd3;
        RAM_1[157] = -16'd6;
        RAM_2[157] = 16'd15;
        RAM_3[157] = -16'd16;
        RAM_0[158] = -16'd20;
        RAM_1[158] = -16'd6;
        RAM_2[158] = -16'd7;
        RAM_3[158] = -16'd5;
        RAM_0[159] = -16'd11;
        RAM_1[159] = 16'd0;
        RAM_2[159] = 16'd0;
        RAM_3[159] = 16'd0;
        RAM_0[160] = -16'd6;
        RAM_1[160] = 16'd6;
        RAM_2[160] = -16'd3;
        RAM_3[160] = -16'd19;
        RAM_0[161] = -16'd1;
        RAM_1[161] = 16'd12;
        RAM_2[161] = 16'd16;
        RAM_3[161] = 16'd6;
        RAM_0[162] = -16'd3;
        RAM_1[162] = -16'd5;
        RAM_2[162] = -16'd5;
        RAM_3[162] = -16'd5;
        RAM_0[163] = -16'd2;
        RAM_1[163] = 16'd1;
        RAM_2[163] = 16'd3;
        RAM_3[163] = 16'd12;
        RAM_0[164] = -16'd6;
        RAM_1[164] = 16'd0;
        RAM_2[164] = 16'd0;
        RAM_3[164] = 16'd0;
        RAM_0[165] = -16'd1;
        RAM_1[165] = -16'd22;
        RAM_2[165] = -16'd2;
        RAM_3[165] = 16'd5;
        RAM_0[166] = 16'd1;
        RAM_1[166] = -16'd2;
        RAM_2[166] = -16'd7;
        RAM_3[166] = 16'd12;
        RAM_0[167] = -16'd3;
        RAM_1[167] = -16'd6;
        RAM_2[167] = -16'd1;
        RAM_3[167] = 16'd7;
        RAM_0[168] = -16'd10;
        RAM_1[168] = -16'd6;
        RAM_2[168] = -16'd1;
        RAM_3[168] = 16'd17;
        RAM_0[169] = 16'd8;
        RAM_1[169] = -16'd13;
        RAM_2[169] = -16'd5;
        RAM_3[169] = -16'd4;
        RAM_0[170] = -16'd9;
        RAM_1[170] = 16'd0;
        RAM_2[170] = 16'd0;
        RAM_3[170] = 16'd0;
        RAM_0[171] = 16'd1;
        RAM_1[171] = -16'd4;
        RAM_2[171] = -16'd5;
        RAM_3[171] = -16'd13;
        RAM_0[172] = -16'd16;
        RAM_1[172] = 16'd0;
        RAM_2[172] = 16'd0;
        RAM_3[172] = 16'd0;
        RAM_0[173] = -16'd19;
        RAM_1[173] = 16'd0;
        RAM_2[173] = -16'd1;
        RAM_3[173] = 16'd13;
        RAM_0[174] = -16'd10;
        RAM_1[174] = 16'd0;
        RAM_2[174] = 16'd0;
        RAM_3[174] = 16'd0;
        RAM_0[175] = -16'd4;
        RAM_1[175] = 16'd0;
        RAM_2[175] = 16'd0;
        RAM_3[175] = 16'd0;
        RAM_0[176] = -16'd29;
        RAM_1[176] = -16'd3;
        RAM_2[176] = 16'd3;
        RAM_3[176] = 16'd6;
        RAM_0[177] = 16'd5;
        RAM_1[177] = -16'd4;
        RAM_2[177] = 16'd4;
        RAM_3[177] = -16'd6;
        RAM_0[178] = -16'd1;
        RAM_1[178] = 16'd9;
        RAM_2[178] = 16'd1;
        RAM_3[178] = 16'd6;
        RAM_0[179] = 16'd0;
        RAM_1[179] = -16'd2;
        RAM_2[179] = -16'd7;
        RAM_3[179] = 16'd21;
        RAM_0[180] = 16'd1;
        RAM_1[180] = -16'd14;
        RAM_2[180] = -16'd27;
        RAM_3[180] = 16'd2;
        RAM_0[181] = 16'd7;
        RAM_1[181] = -16'd2;
        RAM_2[181] = -16'd2;
        RAM_3[181] = 16'd6;
        RAM_0[182] = 16'd4;
        RAM_1[182] = 16'd14;
        RAM_2[182] = 16'd20;
        RAM_3[182] = -16'd5;
        RAM_0[183] = -16'd5;
        RAM_1[183] = 16'd5;
        RAM_2[183] = 16'd4;
        RAM_3[183] = 16'd19;
        RAM_0[184] = 16'd1;
        RAM_1[184] = -16'd10;
        RAM_2[184] = -16'd14;
        RAM_3[184] = -16'd20;
        RAM_0[185] = 16'd8;
        RAM_1[185] = -16'd21;
        RAM_2[185] = -16'd15;
        RAM_3[185] = -16'd3;
        RAM_0[186] = 16'd6;
        RAM_1[186] = -16'd24;
        RAM_2[186] = -16'd11;
        RAM_3[186] = 16'd3;
        RAM_0[187] = 16'd0;
        RAM_1[187] = -16'd2;
        RAM_2[187] = -16'd1;
        RAM_3[187] = 16'd11;
        RAM_0[188] = 16'd2;
        RAM_1[188] = -16'd10;
        RAM_2[188] = 16'd6;
        RAM_3[188] = -16'd6;
        RAM_0[189] = -16'd3;
        RAM_1[189] = 16'd10;
        RAM_2[189] = 16'd1;
        RAM_3[189] = 16'd3;
        RAM_0[190] = -16'd20;
        RAM_1[190] = -16'd9;
        RAM_2[190] = -16'd1;
        RAM_3[190] = -16'd6;
        RAM_0[191] = -16'd11;
        RAM_1[191] = 16'd0;
        RAM_2[191] = 16'd0;
        RAM_3[191] = 16'd0;
        RAM_0[192] = -16'd6;
        RAM_1[192] = 16'd2;
        RAM_2[192] = -16'd6;
        RAM_3[192] = 16'd20;
        RAM_0[193] = -16'd1;
        RAM_1[193] = -16'd4;
        RAM_2[193] = -16'd2;
        RAM_3[193] = -16'd16;
        RAM_0[194] = -16'd3;
        RAM_1[194] = 16'd6;
        RAM_2[194] = 16'd4;
        RAM_3[194] = -16'd20;
        RAM_0[195] = -16'd2;
        RAM_1[195] = -16'd14;
        RAM_2[195] = -16'd14;
        RAM_3[195] = -16'd1;
        RAM_0[196] = -16'd6;
        RAM_1[196] = 16'd0;
        RAM_2[196] = 16'd0;
        RAM_3[196] = 16'd0;
        RAM_0[197] = -16'd1;
        RAM_1[197] = -16'd2;
        RAM_2[197] = -16'd4;
        RAM_3[197] = -16'd6;
        RAM_0[198] = 16'd1;
        RAM_1[198] = -16'd10;
        RAM_2[198] = 16'd0;
        RAM_3[198] = 16'd9;
        RAM_0[199] = -16'd3;
        RAM_1[199] = 16'd7;
        RAM_2[199] = 16'd5;
        RAM_3[199] = -16'd9;
        RAM_0[200] = -16'd10;
        RAM_1[200] = -16'd16;
        RAM_2[200] = -16'd5;
        RAM_3[200] = 16'd19;
        RAM_0[201] = 16'd8;
        RAM_1[201] = -16'd17;
        RAM_2[201] = -16'd5;
        RAM_3[201] = 16'd5;
        RAM_0[202] = -16'd9;
        RAM_1[202] = 16'd0;
        RAM_2[202] = 16'd0;
        RAM_3[202] = 16'd0;
        RAM_0[203] = 16'd1;
        RAM_1[203] = -16'd4;
        RAM_2[203] = -16'd4;
        RAM_3[203] = 16'd16;
        RAM_0[204] = -16'd16;
        RAM_1[204] = 16'd0;
        RAM_2[204] = 16'd0;
        RAM_3[204] = 16'd0;
        RAM_0[205] = -16'd19;
        RAM_1[205] = -16'd9;
        RAM_2[205] = 16'd14;
        RAM_3[205] = -16'd3;
        RAM_0[206] = -16'd10;
        RAM_1[206] = 16'd0;
        RAM_2[206] = 16'd0;
        RAM_3[206] = 16'd0;
        RAM_0[207] = -16'd4;
        RAM_1[207] = 16'd0;
        RAM_2[207] = 16'd0;
        RAM_3[207] = 16'd0;
        RAM_0[208] = -16'd29;
        RAM_1[208] = 16'd8;
        RAM_2[208] = 16'd4;
        RAM_3[208] = 16'd0;
        RAM_0[209] = 16'd5;
        RAM_1[209] = -16'd7;
        RAM_2[209] = 16'd0;
        RAM_3[209] = 16'd14;
        RAM_0[210] = -16'd1;
        RAM_1[210] = -16'd3;
        RAM_2[210] = -16'd9;
        RAM_3[210] = -16'd7;
        RAM_0[211] = 16'd0;
        RAM_1[211] = -16'd12;
        RAM_2[211] = -16'd8;
        RAM_3[211] = 16'd11;
        RAM_0[212] = 16'd1;
        RAM_1[212] = 16'd1;
        RAM_2[212] = 16'd4;
        RAM_3[212] = -16'd14;
        RAM_0[213] = 16'd7;
        RAM_1[213] = -16'd15;
        RAM_2[213] = 16'd5;
        RAM_3[213] = 16'd4;
        RAM_0[214] = 16'd4;
        RAM_1[214] = -16'd2;
        RAM_2[214] = -16'd4;
        RAM_3[214] = -16'd7;
        RAM_0[215] = -16'd5;
        RAM_1[215] = -16'd5;
        RAM_2[215] = 16'd4;
        RAM_3[215] = 16'd24;
        RAM_0[216] = 16'd1;
        RAM_1[216] = 16'd2;
        RAM_2[216] = -16'd7;
        RAM_3[216] = 16'd15;
        RAM_0[217] = 16'd8;
        RAM_1[217] = -16'd26;
        RAM_2[217] = -16'd20;
        RAM_3[217] = 16'd11;
        RAM_0[218] = 16'd6;
        RAM_1[218] = -16'd22;
        RAM_2[218] = -16'd11;
        RAM_3[218] = 16'd2;
        RAM_0[219] = 16'd0;
        RAM_1[219] = -16'd11;
        RAM_2[219] = -16'd2;
        RAM_3[219] = 16'd5;
        RAM_0[220] = 16'd2;
        RAM_1[220] = -16'd24;
        RAM_2[220] = -16'd13;
        RAM_3[220] = 16'd2;
        RAM_0[221] = -16'd3;
        RAM_1[221] = -16'd6;
        RAM_2[221] = -16'd6;
        RAM_3[221] = 16'd13;
        RAM_0[222] = -16'd20;
        RAM_1[222] = 16'd6;
        RAM_2[222] = -16'd2;
        RAM_3[222] = 16'd1;
        RAM_0[223] = -16'd11;
        RAM_1[223] = 16'd0;
        RAM_2[223] = 16'd0;
        RAM_3[223] = 16'd0;
        RAM_0[224] = -16'd6;
        RAM_1[224] = 16'd1;
        RAM_2[224] = -16'd3;
        RAM_3[224] = -16'd3;
        RAM_0[225] = -16'd1;
        RAM_1[225] = 16'd0;
        RAM_2[225] = 16'd1;
        RAM_3[225] = 16'd2;
        RAM_0[226] = -16'd3;
        RAM_1[226] = 16'd0;
        RAM_2[226] = -16'd1;
        RAM_3[226] = 16'd0;
        RAM_0[227] = -16'd2;
        RAM_1[227] = 16'd0;
        RAM_2[227] = 16'd0;
        RAM_3[227] = 16'd1;
        RAM_0[228] = -16'd6;
        RAM_1[228] = 16'd0;
        RAM_2[228] = 16'd0;
        RAM_3[228] = 16'd0;
        RAM_0[229] = -16'd1;
        RAM_1[229] = -16'd1;
        RAM_2[229] = -16'd1;
        RAM_3[229] = -16'd5;
        RAM_0[230] = 16'd1;
        RAM_1[230] = 16'd0;
        RAM_2[230] = -16'd6;
        RAM_3[230] = 16'd4;
        RAM_0[231] = -16'd3;
        RAM_1[231] = 16'd1;
        RAM_2[231] = -16'd2;
        RAM_3[231] = 16'd9;
        RAM_0[232] = -16'd10;
        RAM_1[232] = -16'd12;
        RAM_2[232] = -16'd1;
        RAM_3[232] = -16'd2;
        RAM_0[233] = 16'd8;
        RAM_1[233] = -16'd16;
        RAM_2[233] = -16'd7;
        RAM_3[233] = -16'd2;
        RAM_0[234] = -16'd9;
        RAM_1[234] = 16'd0;
        RAM_2[234] = 16'd0;
        RAM_3[234] = 16'd0;
        RAM_0[235] = 16'd1;
        RAM_1[235] = 16'd0;
        RAM_2[235] = -16'd1;
        RAM_3[235] = 16'd4;
        RAM_0[236] = -16'd16;
        RAM_1[236] = 16'd0;
        RAM_2[236] = 16'd0;
        RAM_3[236] = 16'd0;
        RAM_0[237] = -16'd19;
        RAM_1[237] = -16'd5;
        RAM_2[237] = 16'd0;
        RAM_3[237] = 16'd0;
        RAM_0[238] = -16'd10;
        RAM_1[238] = 16'd0;
        RAM_2[238] = 16'd0;
        RAM_3[238] = 16'd0;
        RAM_0[239] = -16'd4;
        RAM_1[239] = 16'd0;
        RAM_2[239] = 16'd0;
        RAM_3[239] = 16'd0;
        RAM_0[240] = -16'd29;
        RAM_1[240] = -16'd2;
        RAM_2[240] = 16'd0;
        RAM_3[240] = 16'd0;
        RAM_0[241] = 16'd5;
        RAM_1[241] = -16'd15;
        RAM_2[241] = -16'd8;
        RAM_3[241] = -16'd2;
        RAM_0[242] = -16'd1;
        RAM_1[242] = 16'd0;
        RAM_2[242] = 16'd0;
        RAM_3[242] = 16'd0;
        RAM_0[243] = 16'd0;
        RAM_1[243] = -16'd6;
        RAM_2[243] = 16'd1;
        RAM_3[243] = 16'd0;
        RAM_0[244] = 16'd1;
        RAM_1[244] = 16'd0;
        RAM_2[244] = 16'd0;
        RAM_3[244] = -16'd5;
        RAM_0[245] = 16'd7;
        RAM_1[245] = -16'd27;
        RAM_2[245] = -16'd2;
        RAM_3[245] = -16'd1;
        RAM_0[246] = 16'd4;
        RAM_1[246] = 16'd0;
        RAM_2[246] = -16'd2;
        RAM_3[246] = 16'd2;
        RAM_0[247] = -16'd5;
        RAM_1[247] = -16'd13;
        RAM_2[247] = -16'd13;
        RAM_3[247] = -16'd5;
        RAM_0[248] = 16'd1;
        RAM_1[248] = 16'd0;
        RAM_2[248] = 16'd0;
        RAM_3[248] = -16'd4;
        RAM_0[249] = 16'd8;
        RAM_1[249] = -16'd17;
        RAM_2[249] = -16'd6;
        RAM_3[249] = -16'd6;
        RAM_0[250] = 16'd6;
        RAM_1[250] = -16'd20;
        RAM_2[250] = -16'd3;
        RAM_3[250] = -16'd2;
        RAM_0[251] = 16'd0;
        RAM_1[251] = -16'd8;
        RAM_2[251] = -16'd4;
        RAM_3[251] = 16'd2;
        RAM_0[252] = 16'd2;
        RAM_1[252] = -16'd19;
        RAM_2[252] = -16'd6;
        RAM_3[252] = 16'd0;
        RAM_0[253] = -16'd3;
        RAM_1[253] = 16'd0;
        RAM_2[253] = -16'd3;
        RAM_3[253] = -16'd10;
        RAM_0[254] = -16'd20;
        RAM_1[254] = 16'd12;
        RAM_2[254] = 16'd7;
        RAM_3[254] = 16'd2;
        RAM_0[255] = -16'd11;
        RAM_1[255] = 16'd0;
        RAM_2[255] = 16'd0;
        RAM_3[255] = 16'd0;
        RAM_0[256] = -16'd6;
        RAM_1[256] = 16'd0;
        RAM_2[256] = -16'd20;
        RAM_3[256] = -16'd10;
        RAM_0[257] = -16'd1;
        RAM_1[257] = -16'd2;
        RAM_2[257] = -16'd9;
        RAM_3[257] = -16'd17;
        RAM_0[258] = -16'd3;
        RAM_1[258] = -16'd1;
        RAM_2[258] = -16'd2;
        RAM_3[258] = -16'd7;
        RAM_0[259] = -16'd2;
        RAM_1[259] = -16'd6;
        RAM_2[259] = 16'd7;
        RAM_3[259] = -16'd20;
        RAM_0[260] = -16'd6;
        RAM_1[260] = 16'd0;
        RAM_2[260] = 16'd0;
        RAM_3[260] = 16'd0;
        RAM_0[261] = -16'd1;
        RAM_1[261] = 16'd6;
        RAM_2[261] = -16'd2;
        RAM_3[261] = -16'd3;
        RAM_0[262] = 16'd1;
        RAM_1[262] = 16'd0;
        RAM_2[262] = -16'd22;
        RAM_3[262] = -16'd4;
        RAM_0[263] = -16'd3;
        RAM_1[263] = -16'd1;
        RAM_2[263] = -16'd5;
        RAM_3[263] = -16'd7;
        RAM_0[264] = -16'd10;
        RAM_1[264] = -16'd11;
        RAM_2[264] = -16'd2;
        RAM_3[264] = 16'd7;
        RAM_0[265] = 16'd8;
        RAM_1[265] = 16'd0;
        RAM_2[265] = 16'd7;
        RAM_3[265] = -16'd6;
        RAM_0[266] = -16'd9;
        RAM_1[266] = 16'd0;
        RAM_2[266] = 16'd0;
        RAM_3[266] = 16'd0;
        RAM_0[267] = 16'd1;
        RAM_1[267] = 16'd1;
        RAM_2[267] = -16'd26;
        RAM_3[267] = -16'd3;
        RAM_0[268] = -16'd16;
        RAM_1[268] = 16'd0;
        RAM_2[268] = 16'd0;
        RAM_3[268] = 16'd0;
        RAM_0[269] = -16'd19;
        RAM_1[269] = 16'd11;
        RAM_2[269] = 16'd10;
        RAM_3[269] = -16'd4;
        RAM_0[270] = -16'd10;
        RAM_1[270] = 16'd0;
        RAM_2[270] = 16'd0;
        RAM_3[270] = 16'd0;
        RAM_0[271] = -16'd4;
        RAM_1[271] = 16'd0;
        RAM_2[271] = 16'd0;
        RAM_3[271] = 16'd0;
        RAM_0[272] = -16'd29;
        RAM_1[272] = 16'd14;
        RAM_2[272] = 16'd9;
        RAM_3[272] = 16'd3;
        RAM_0[273] = 16'd5;
        RAM_1[273] = 16'd0;
        RAM_2[273] = -16'd11;
        RAM_3[273] = 16'd4;
        RAM_0[274] = -16'd1;
        RAM_1[274] = -16'd2;
        RAM_2[274] = -16'd31;
        RAM_3[274] = 16'd0;
        RAM_0[275] = 16'd0;
        RAM_1[275] = -16'd5;
        RAM_2[275] = -16'd7;
        RAM_3[275] = 16'd1;
        RAM_0[276] = 16'd1;
        RAM_1[276] = -16'd21;
        RAM_2[276] = -16'd16;
        RAM_3[276] = 16'd4;
        RAM_0[277] = 16'd7;
        RAM_1[277] = -16'd2;
        RAM_2[277] = 16'd9;
        RAM_3[277] = -16'd6;
        RAM_0[278] = 16'd4;
        RAM_1[278] = 16'd0;
        RAM_2[278] = -16'd7;
        RAM_3[278] = -16'd16;
        RAM_0[279] = -16'd5;
        RAM_1[279] = -16'd1;
        RAM_2[279] = -16'd6;
        RAM_3[279] = 16'd9;
        RAM_0[280] = 16'd1;
        RAM_1[280] = -16'd3;
        RAM_2[280] = -16'd4;
        RAM_3[280] = -16'd2;
        RAM_0[281] = 16'd8;
        RAM_1[281] = 16'd0;
        RAM_2[281] = 16'd1;
        RAM_3[281] = -16'd7;
        RAM_0[282] = 16'd6;
        RAM_1[282] = 16'd0;
        RAM_2[282] = 16'd8;
        RAM_3[282] = -16'd15;
        RAM_0[283] = 16'd0;
        RAM_1[283] = 16'd1;
        RAM_2[283] = -16'd16;
        RAM_3[283] = 16'd13;
        RAM_0[284] = 16'd2;
        RAM_1[284] = 16'd0;
        RAM_2[284] = -16'd13;
        RAM_3[284] = -16'd1;
        RAM_0[285] = -16'd3;
        RAM_1[285] = -16'd3;
        RAM_2[285] = -16'd21;
        RAM_3[285] = -16'd7;
        RAM_0[286] = -16'd20;
        RAM_1[286] = -16'd6;
        RAM_2[286] = -16'd1;
        RAM_3[286] = 16'd1;
        RAM_0[287] = -16'd11;
        RAM_1[287] = 16'd0;
        RAM_2[287] = 16'd0;
        RAM_3[287] = 16'd0;
        RAM_0[288] = -16'd6;
        RAM_1[288] = 16'd5;
        RAM_2[288] = -16'd19;
        RAM_3[288] = -16'd15;
        RAM_0[289] = -16'd1;
        RAM_1[289] = 16'd3;
        RAM_2[289] = -16'd2;
        RAM_3[289] = -16'd31;
        RAM_0[290] = -16'd3;
        RAM_1[290] = 16'd15;
        RAM_2[290] = 16'd4;
        RAM_3[290] = -16'd22;
        RAM_0[291] = -16'd2;
        RAM_1[291] = 16'd9;
        RAM_2[291] = -16'd10;
        RAM_3[291] = -16'd4;
        RAM_0[292] = -16'd6;
        RAM_1[292] = 16'd0;
        RAM_2[292] = 16'd0;
        RAM_3[292] = 16'd0;
        RAM_0[293] = -16'd1;
        RAM_1[293] = 16'd16;
        RAM_2[293] = -16'd7;
        RAM_3[293] = -16'd1;
        RAM_0[294] = 16'd1;
        RAM_1[294] = 16'd11;
        RAM_2[294] = -16'd29;
        RAM_3[294] = -16'd39;
        RAM_0[295] = -16'd3;
        RAM_1[295] = 16'd11;
        RAM_2[295] = 16'd1;
        RAM_3[295] = -16'd24;
        RAM_0[296] = -16'd10;
        RAM_1[296] = -16'd1;
        RAM_2[296] = -16'd8;
        RAM_3[296] = -16'd10;
        RAM_0[297] = 16'd8;
        RAM_1[297] = 16'd10;
        RAM_2[297] = -16'd8;
        RAM_3[297] = -16'd9;
        RAM_0[298] = -16'd9;
        RAM_1[298] = 16'd0;
        RAM_2[298] = 16'd0;
        RAM_3[298] = 16'd0;
        RAM_0[299] = 16'd1;
        RAM_1[299] = 16'd9;
        RAM_2[299] = -16'd14;
        RAM_3[299] = -16'd17;
        RAM_0[300] = -16'd16;
        RAM_1[300] = 16'd0;
        RAM_2[300] = 16'd0;
        RAM_3[300] = 16'd0;
        RAM_0[301] = -16'd19;
        RAM_1[301] = -16'd5;
        RAM_2[301] = 16'd0;
        RAM_3[301] = 16'd15;
        RAM_0[302] = -16'd10;
        RAM_1[302] = 16'd0;
        RAM_2[302] = 16'd0;
        RAM_3[302] = 16'd0;
        RAM_0[303] = -16'd4;
        RAM_1[303] = 16'd0;
        RAM_2[303] = 16'd0;
        RAM_3[303] = 16'd0;
        RAM_0[304] = -16'd29;
        RAM_1[304] = -16'd2;
        RAM_2[304] = 16'd2;
        RAM_3[304] = -16'd14;
        RAM_0[305] = 16'd5;
        RAM_1[305] = 16'd5;
        RAM_2[305] = -16'd3;
        RAM_3[305] = -16'd14;
        RAM_0[306] = -16'd1;
        RAM_1[306] = 16'd8;
        RAM_2[306] = -16'd11;
        RAM_3[306] = -16'd9;
        RAM_0[307] = 16'd0;
        RAM_1[307] = 16'd3;
        RAM_2[307] = -16'd3;
        RAM_3[307] = -16'd18;
        RAM_0[308] = 16'd1;
        RAM_1[308] = 16'd6;
        RAM_2[308] = -16'd2;
        RAM_3[308] = -16'd45;
        RAM_0[309] = 16'd7;
        RAM_1[309] = 16'd12;
        RAM_2[309] = 16'd3;
        RAM_3[309] = -16'd22;
        RAM_0[310] = 16'd4;
        RAM_1[310] = 16'd3;
        RAM_2[310] = -16'd18;
        RAM_3[310] = -16'd23;
        RAM_0[311] = -16'd5;
        RAM_1[311] = 16'd4;
        RAM_2[311] = -16'd6;
        RAM_3[311] = -16'd13;
        RAM_0[312] = 16'd1;
        RAM_1[312] = 16'd8;
        RAM_2[312] = -16'd7;
        RAM_3[312] = 16'd0;
        RAM_0[313] = 16'd8;
        RAM_1[313] = -16'd5;
        RAM_2[313] = -16'd6;
        RAM_3[313] = -16'd17;
        RAM_0[314] = 16'd6;
        RAM_1[314] = 16'd7;
        RAM_2[314] = -16'd7;
        RAM_3[314] = -16'd11;
        RAM_0[315] = 16'd0;
        RAM_1[315] = -16'd7;
        RAM_2[315] = -16'd4;
        RAM_3[315] = -16'd25;
        RAM_0[316] = 16'd2;
        RAM_1[316] = 16'd2;
        RAM_2[316] = -16'd16;
        RAM_3[316] = 16'd1;
        RAM_0[317] = -16'd3;
        RAM_1[317] = 16'd7;
        RAM_2[317] = -16'd28;
        RAM_3[317] = -16'd31;
        RAM_0[318] = -16'd20;
        RAM_1[318] = -16'd7;
        RAM_2[318] = 16'd1;
        RAM_3[318] = -16'd9;
        RAM_0[319] = -16'd11;
        RAM_1[319] = 16'd0;
        RAM_2[319] = 16'd0;
        RAM_3[319] = 16'd0;
        RAM_0[320] = -16'd6;
        RAM_1[320] = -16'd3;
        RAM_2[320] = 16'd0;
        RAM_3[320] = 16'd1;
        RAM_0[321] = -16'd1;
        RAM_1[321] = -16'd8;
        RAM_2[321] = -16'd6;
        RAM_3[321] = 16'd4;
        RAM_0[322] = -16'd3;
        RAM_1[322] = -16'd4;
        RAM_2[322] = -16'd6;
        RAM_3[322] = 16'd0;
        RAM_0[323] = -16'd2;
        RAM_1[323] = 16'd5;
        RAM_2[323] = -16'd2;
        RAM_3[323] = -16'd2;
        RAM_0[324] = -16'd6;
        RAM_1[324] = 16'd0;
        RAM_2[324] = 16'd0;
        RAM_3[324] = 16'd0;
        RAM_0[325] = -16'd1;
        RAM_1[325] = 16'd10;
        RAM_2[325] = -16'd20;
        RAM_3[325] = -16'd26;
        RAM_0[326] = 16'd1;
        RAM_1[326] = -16'd2;
        RAM_2[326] = -16'd10;
        RAM_3[326] = 16'd8;
        RAM_0[327] = -16'd3;
        RAM_1[327] = -16'd5;
        RAM_2[327] = -16'd6;
        RAM_3[327] = 16'd7;
        RAM_0[328] = -16'd10;
        RAM_1[328] = 16'd3;
        RAM_2[328] = -16'd7;
        RAM_3[328] = 16'd0;
        RAM_0[329] = 16'd8;
        RAM_1[329] = -16'd1;
        RAM_2[329] = -16'd8;
        RAM_3[329] = -16'd18;
        RAM_0[330] = -16'd9;
        RAM_1[330] = 16'd0;
        RAM_2[330] = 16'd0;
        RAM_3[330] = 16'd0;
        RAM_0[331] = 16'd1;
        RAM_1[331] = 16'd2;
        RAM_2[331] = -16'd2;
        RAM_3[331] = -16'd3;
        RAM_0[332] = -16'd16;
        RAM_1[332] = 16'd0;
        RAM_2[332] = 16'd0;
        RAM_3[332] = 16'd0;
        RAM_0[333] = -16'd19;
        RAM_1[333] = 16'd0;
        RAM_2[333] = 16'd0;
        RAM_3[333] = 16'd8;
        RAM_0[334] = -16'd10;
        RAM_1[334] = 16'd0;
        RAM_2[334] = 16'd0;
        RAM_3[334] = 16'd0;
        RAM_0[335] = -16'd4;
        RAM_1[335] = 16'd0;
        RAM_2[335] = 16'd0;
        RAM_3[335] = 16'd0;
        RAM_0[336] = -16'd29;
        RAM_1[336] = -16'd6;
        RAM_2[336] = -16'd5;
        RAM_3[336] = 16'd3;
        RAM_0[337] = 16'd5;
        RAM_1[337] = -16'd6;
        RAM_2[337] = -16'd7;
        RAM_3[337] = -16'd9;
        RAM_0[338] = -16'd1;
        RAM_1[338] = 16'd1;
        RAM_2[338] = 16'd0;
        RAM_3[338] = -16'd6;
        RAM_0[339] = 16'd0;
        RAM_1[339] = -16'd9;
        RAM_2[339] = -16'd10;
        RAM_3[339] = 16'd2;
        RAM_0[340] = 16'd1;
        RAM_1[340] = 16'd6;
        RAM_2[340] = -16'd11;
        RAM_3[340] = 16'd6;
        RAM_0[341] = 16'd7;
        RAM_1[341] = -16'd9;
        RAM_2[341] = -16'd17;
        RAM_3[341] = -16'd10;
        RAM_0[342] = 16'd4;
        RAM_1[342] = -16'd16;
        RAM_2[342] = -16'd13;
        RAM_3[342] = 16'd6;
        RAM_0[343] = -16'd5;
        RAM_1[343] = -16'd9;
        RAM_2[343] = -16'd16;
        RAM_3[343] = 16'd0;
        RAM_0[344] = 16'd1;
        RAM_1[344] = 16'd0;
        RAM_2[344] = 16'd2;
        RAM_3[344] = -16'd1;
        RAM_0[345] = 16'd8;
        RAM_1[345] = -16'd1;
        RAM_2[345] = -16'd2;
        RAM_3[345] = -16'd26;
        RAM_0[346] = 16'd6;
        RAM_1[346] = 16'd0;
        RAM_2[346] = -16'd9;
        RAM_3[346] = -16'd30;
        RAM_0[347] = 16'd0;
        RAM_1[347] = -16'd22;
        RAM_2[347] = -16'd21;
        RAM_3[347] = 16'd4;
        RAM_0[348] = 16'd2;
        RAM_1[348] = 16'd3;
        RAM_2[348] = -16'd5;
        RAM_3[348] = -16'd15;
        RAM_0[349] = -16'd3;
        RAM_1[349] = 16'd3;
        RAM_2[349] = -16'd7;
        RAM_3[349] = 16'd1;
        RAM_0[350] = -16'd20;
        RAM_1[350] = 16'd19;
        RAM_2[350] = 16'd3;
        RAM_3[350] = 16'd5;
        RAM_0[351] = -16'd11;
        RAM_1[351] = 16'd0;
        RAM_2[351] = 16'd0;
        RAM_3[351] = 16'd0;
        RAM_0[352] = -16'd6;
        RAM_1[352] = -16'd26;
        RAM_2[352] = -16'd17;
        RAM_3[352] = -16'd11;
        RAM_0[353] = -16'd1;
        RAM_1[353] = -16'd37;
        RAM_2[353] = -16'd21;
        RAM_3[353] = -16'd19;
        RAM_0[354] = -16'd3;
        RAM_1[354] = -16'd35;
        RAM_2[354] = -16'd28;
        RAM_3[354] = -16'd31;
        RAM_0[355] = -16'd2;
        RAM_1[355] = -16'd33;
        RAM_2[355] = -16'd21;
        RAM_3[355] = -16'd3;
        RAM_0[356] = -16'd6;
        RAM_1[356] = 16'd0;
        RAM_2[356] = 16'd0;
        RAM_3[356] = 16'd0;
        RAM_0[357] = -16'd1;
        RAM_1[357] = 16'd1;
        RAM_2[357] = -16'd9;
        RAM_3[357] = 16'd5;
        RAM_0[358] = 16'd1;
        RAM_1[358] = -16'd30;
        RAM_2[358] = -16'd25;
        RAM_3[358] = -16'd7;
        RAM_0[359] = -16'd3;
        RAM_1[359] = -16'd35;
        RAM_2[359] = -16'd26;
        RAM_3[359] = -16'd26;
        RAM_0[360] = -16'd10;
        RAM_1[360] = 16'd10;
        RAM_2[360] = -16'd3;
        RAM_3[360] = -16'd4;
        RAM_0[361] = 16'd8;
        RAM_1[361] = -16'd1;
        RAM_2[361] = 16'd6;
        RAM_3[361] = -16'd5;
        RAM_0[362] = -16'd9;
        RAM_1[362] = 16'd0;
        RAM_2[362] = 16'd0;
        RAM_3[362] = 16'd0;
        RAM_0[363] = 16'd1;
        RAM_1[363] = -16'd28;
        RAM_2[363] = -16'd28;
        RAM_3[363] = -16'd13;
        RAM_0[364] = -16'd16;
        RAM_1[364] = 16'd0;
        RAM_2[364] = 16'd0;
        RAM_3[364] = 16'd0;
        RAM_0[365] = -16'd19;
        RAM_1[365] = 16'd11;
        RAM_2[365] = -16'd18;
        RAM_3[365] = 16'd2;
        RAM_0[366] = -16'd10;
        RAM_1[366] = 16'd0;
        RAM_2[366] = 16'd0;
        RAM_3[366] = 16'd0;
        RAM_0[367] = -16'd4;
        RAM_1[367] = 16'd0;
        RAM_2[367] = 16'd0;
        RAM_3[367] = 16'd0;
        RAM_0[368] = -16'd29;
        RAM_1[368] = 16'd2;
        RAM_2[368] = -16'd3;
        RAM_3[368] = 16'd0;
        RAM_0[369] = 16'd5;
        RAM_1[369] = 16'd3;
        RAM_2[369] = 16'd2;
        RAM_3[369] = -16'd5;
        RAM_0[370] = -16'd1;
        RAM_1[370] = -16'd25;
        RAM_2[370] = -16'd27;
        RAM_3[370] = -16'd10;
        RAM_0[371] = 16'd0;
        RAM_1[371] = 16'd6;
        RAM_2[371] = 16'd1;
        RAM_3[371] = 16'd0;
        RAM_0[372] = 16'd1;
        RAM_1[372] = -16'd26;
        RAM_2[372] = -16'd36;
        RAM_3[372] = -16'd19;
        RAM_0[373] = 16'd7;
        RAM_1[373] = 16'd3;
        RAM_2[373] = -16'd4;
        RAM_3[373] = 16'd1;
        RAM_0[374] = 16'd4;
        RAM_1[374] = -16'd31;
        RAM_2[374] = -16'd31;
        RAM_3[374] = -16'd20;
        RAM_0[375] = -16'd5;
        RAM_1[375] = 16'd13;
        RAM_2[375] = -16'd3;
        RAM_3[375] = -16'd19;
        RAM_0[376] = 16'd1;
        RAM_1[376] = -16'd36;
        RAM_2[376] = -16'd29;
        RAM_3[376] = -16'd4;
        RAM_0[377] = 16'd8;
        RAM_1[377] = -16'd3;
        RAM_2[377] = 16'd7;
        RAM_3[377] = 16'd5;
        RAM_0[378] = 16'd6;
        RAM_1[378] = -16'd6;
        RAM_2[378] = 16'd12;
        RAM_3[378] = 16'd0;
        RAM_0[379] = 16'd0;
        RAM_1[379] = 16'd17;
        RAM_2[379] = -16'd3;
        RAM_3[379] = -16'd9;
        RAM_0[380] = 16'd2;
        RAM_1[380] = -16'd4;
        RAM_2[380] = 16'd8;
        RAM_3[380] = -16'd5;
        RAM_0[381] = -16'd3;
        RAM_1[381] = -16'd28;
        RAM_2[381] = -16'd21;
        RAM_3[381] = -16'd6;
        RAM_0[382] = -16'd20;
        RAM_1[382] = -16'd1;
        RAM_2[382] = 16'd4;
        RAM_3[382] = -16'd10;
        RAM_0[383] = -16'd11;
        RAM_1[383] = 16'd0;
        RAM_2[383] = 16'd0;
        RAM_3[383] = 16'd0;
        RAM_0[384] = -16'd6;
        RAM_1[384] = -16'd11;
        RAM_2[384] = -16'd10;
        RAM_3[384] = 16'd9;
        RAM_0[385] = -16'd1;
        RAM_1[385] = 16'd4;
        RAM_2[385] = -16'd4;
        RAM_3[385] = 16'd1;
        RAM_0[386] = -16'd3;
        RAM_1[386] = -16'd3;
        RAM_2[386] = -16'd7;
        RAM_3[386] = 16'd1;
        RAM_0[387] = -16'd2;
        RAM_1[387] = -16'd10;
        RAM_2[387] = 16'd14;
        RAM_3[387] = -16'd4;
        RAM_0[388] = -16'd6;
        RAM_1[388] = 16'd0;
        RAM_2[388] = 16'd0;
        RAM_3[388] = 16'd0;
        RAM_0[389] = -16'd1;
        RAM_1[389] = -16'd1;
        RAM_2[389] = 16'd0;
        RAM_3[389] = -16'd4;
        RAM_0[390] = 16'd1;
        RAM_1[390] = -16'd14;
        RAM_2[390] = -16'd16;
        RAM_3[390] = 16'd5;
        RAM_0[391] = -16'd3;
        RAM_1[391] = 16'd3;
        RAM_2[391] = -16'd1;
        RAM_3[391] = -16'd2;
        RAM_0[392] = -16'd10;
        RAM_1[392] = 16'd3;
        RAM_2[392] = -16'd7;
        RAM_3[392] = -16'd1;
        RAM_0[393] = 16'd8;
        RAM_1[393] = 16'd13;
        RAM_2[393] = 16'd7;
        RAM_3[393] = 16'd8;
        RAM_0[394] = -16'd9;
        RAM_1[394] = 16'd0;
        RAM_2[394] = 16'd0;
        RAM_3[394] = 16'd0;
        RAM_0[395] = 16'd1;
        RAM_1[395] = -16'd11;
        RAM_2[395] = -16'd16;
        RAM_3[395] = 16'd1;
        RAM_0[396] = -16'd16;
        RAM_1[396] = 16'd0;
        RAM_2[396] = 16'd0;
        RAM_3[396] = 16'd0;
        RAM_0[397] = -16'd19;
        RAM_1[397] = 16'd7;
        RAM_2[397] = -16'd8;
        RAM_3[397] = -16'd1;
        RAM_0[398] = -16'd10;
        RAM_1[398] = 16'd0;
        RAM_2[398] = 16'd0;
        RAM_3[398] = 16'd0;
        RAM_0[399] = -16'd4;
        RAM_1[399] = 16'd0;
        RAM_2[399] = 16'd0;
        RAM_3[399] = 16'd0;
        RAM_0[400] = -16'd29;
        RAM_1[400] = -16'd2;
        RAM_2[400] = 16'd0;
        RAM_3[400] = 16'd0;
        RAM_0[401] = 16'd5;
        RAM_1[401] = 16'd9;
        RAM_2[401] = 16'd4;
        RAM_3[401] = 16'd9;
        RAM_0[402] = -16'd1;
        RAM_1[402] = -16'd9;
        RAM_2[402] = -16'd8;
        RAM_3[402] = 16'd3;
        RAM_0[403] = 16'd0;
        RAM_1[403] = 16'd3;
        RAM_2[403] = -16'd3;
        RAM_3[403] = 16'd4;
        RAM_0[404] = 16'd1;
        RAM_1[404] = -16'd11;
        RAM_2[404] = -16'd11;
        RAM_3[404] = 16'd5;
        RAM_0[405] = 16'd7;
        RAM_1[405] = 16'd17;
        RAM_2[405] = 16'd5;
        RAM_3[405] = 16'd14;
        RAM_0[406] = 16'd4;
        RAM_1[406] = -16'd4;
        RAM_2[406] = -16'd15;
        RAM_3[406] = -16'd5;
        RAM_0[407] = -16'd5;
        RAM_1[407] = 16'd3;
        RAM_2[407] = -16'd3;
        RAM_3[407] = 16'd8;
        RAM_0[408] = 16'd1;
        RAM_1[408] = -16'd9;
        RAM_2[408] = 16'd6;
        RAM_3[408] = 16'd2;
        RAM_0[409] = 16'd8;
        RAM_1[409] = 16'd16;
        RAM_2[409] = 16'd6;
        RAM_3[409] = 16'd11;
        RAM_0[410] = 16'd6;
        RAM_1[410] = 16'd18;
        RAM_2[410] = 16'd5;
        RAM_3[410] = 16'd8;
        RAM_0[411] = 16'd0;
        RAM_1[411] = 16'd0;
        RAM_2[411] = -16'd2;
        RAM_3[411] = 16'd7;
        RAM_0[412] = 16'd2;
        RAM_1[412] = 16'd12;
        RAM_2[412] = 16'd5;
        RAM_3[412] = -16'd1;
        RAM_0[413] = -16'd3;
        RAM_1[413] = -16'd9;
        RAM_2[413] = -16'd7;
        RAM_3[413] = -16'd1;
        RAM_0[414] = -16'd20;
        RAM_1[414] = 16'd1;
        RAM_2[414] = 16'd10;
        RAM_3[414] = 16'd9;
        RAM_0[415] = -16'd11;
        RAM_1[415] = 16'd0;
        RAM_2[415] = 16'd0;
        RAM_3[415] = 16'd0;
        RAM_0[416] = -16'd6;
        RAM_1[416] = -16'd29;
        RAM_2[416] = -16'd3;
        RAM_3[416] = 16'd0;
        RAM_0[417] = -16'd1;
        RAM_1[417] = -16'd26;
        RAM_2[417] = -16'd14;
        RAM_3[417] = -16'd12;
        RAM_0[418] = -16'd3;
        RAM_1[418] = -16'd34;
        RAM_2[418] = -16'd13;
        RAM_3[418] = -16'd10;
        RAM_0[419] = -16'd2;
        RAM_1[419] = -16'd24;
        RAM_2[419] = -16'd8;
        RAM_3[419] = -16'd2;
        RAM_0[420] = -16'd6;
        RAM_1[420] = 16'd0;
        RAM_2[420] = 16'd0;
        RAM_3[420] = 16'd0;
        RAM_0[421] = -16'd1;
        RAM_1[421] = -16'd2;
        RAM_2[421] = -16'd9;
        RAM_3[421] = 16'd10;
        RAM_0[422] = 16'd1;
        RAM_1[422] = -16'd38;
        RAM_2[422] = -16'd14;
        RAM_3[422] = 16'd3;
        RAM_0[423] = -16'd3;
        RAM_1[423] = -16'd27;
        RAM_2[423] = -16'd14;
        RAM_3[423] = -16'd7;
        RAM_0[424] = -16'd10;
        RAM_1[424] = -16'd2;
        RAM_2[424] = -16'd7;
        RAM_3[424] = 16'd1;
        RAM_0[425] = 16'd8;
        RAM_1[425] = 16'd5;
        RAM_2[425] = 16'd0;
        RAM_3[425] = 16'd10;
        RAM_0[426] = -16'd9;
        RAM_1[426] = 16'd0;
        RAM_2[426] = 16'd0;
        RAM_3[426] = 16'd0;
        RAM_0[427] = 16'd1;
        RAM_1[427] = -16'd23;
        RAM_2[427] = -16'd16;
        RAM_3[427] = -16'd20;
        RAM_0[428] = -16'd16;
        RAM_1[428] = 16'd0;
        RAM_2[428] = 16'd0;
        RAM_3[428] = 16'd0;
        RAM_0[429] = -16'd19;
        RAM_1[429] = 16'd5;
        RAM_2[429] = -16'd9;
        RAM_3[429] = -16'd1;
        RAM_0[430] = -16'd10;
        RAM_1[430] = 16'd0;
        RAM_2[430] = 16'd0;
        RAM_3[430] = 16'd0;
        RAM_0[431] = -16'd4;
        RAM_1[431] = 16'd0;
        RAM_2[431] = 16'd0;
        RAM_3[431] = 16'd0;
        RAM_0[432] = -16'd29;
        RAM_1[432] = 16'd9;
        RAM_2[432] = 16'd3;
        RAM_3[432] = 16'd0;
        RAM_0[433] = 16'd5;
        RAM_1[433] = -16'd1;
        RAM_2[433] = -16'd6;
        RAM_3[433] = 16'd9;
        RAM_0[434] = -16'd1;
        RAM_1[434] = -16'd23;
        RAM_2[434] = -16'd17;
        RAM_3[434] = -16'd14;
        RAM_0[435] = 16'd0;
        RAM_1[435] = 16'd0;
        RAM_2[435] = -16'd11;
        RAM_3[435] = 16'd8;
        RAM_0[436] = 16'd1;
        RAM_1[436] = -16'd39;
        RAM_2[436] = -16'd18;
        RAM_3[436] = -16'd8;
        RAM_0[437] = 16'd7;
        RAM_1[437] = 16'd1;
        RAM_2[437] = -16'd4;
        RAM_3[437] = 16'd6;
        RAM_0[438] = 16'd4;
        RAM_1[438] = -16'd24;
        RAM_2[438] = -16'd25;
        RAM_3[438] = -16'd8;
        RAM_0[439] = -16'd5;
        RAM_1[439] = -16'd11;
        RAM_2[439] = -16'd12;
        RAM_3[439] = 16'd2;
        RAM_0[440] = 16'd1;
        RAM_1[440] = -16'd14;
        RAM_2[440] = -16'd2;
        RAM_3[440] = -16'd14;
        RAM_0[441] = 16'd8;
        RAM_1[441] = 16'd9;
        RAM_2[441] = -16'd3;
        RAM_3[441] = 16'd4;
        RAM_0[442] = 16'd6;
        RAM_1[442] = 16'd2;
        RAM_2[442] = 16'd1;
        RAM_3[442] = 16'd3;
        RAM_0[443] = 16'd0;
        RAM_1[443] = -16'd1;
        RAM_2[443] = -16'd3;
        RAM_3[443] = -16'd3;
        RAM_0[444] = 16'd2;
        RAM_1[444] = 16'd3;
        RAM_2[444] = -16'd2;
        RAM_3[444] = -16'd3;
        RAM_0[445] = -16'd3;
        RAM_1[445] = -16'd24;
        RAM_2[445] = -16'd11;
        RAM_3[445] = 16'd1;
        RAM_0[446] = -16'd20;
        RAM_1[446] = 16'd21;
        RAM_2[446] = 16'd4;
        RAM_3[446] = -16'd1;
        RAM_0[447] = -16'd11;
        RAM_1[447] = 16'd0;
        RAM_2[447] = 16'd0;
        RAM_3[447] = 16'd0;
        RAM_0[448] = -16'd6;
        RAM_1[448] = -16'd5;
        RAM_2[448] = -16'd16;
        RAM_3[448] = 16'd6;
        RAM_0[449] = -16'd1;
        RAM_1[449] = 16'd4;
        RAM_2[449] = -16'd10;
        RAM_3[449] = 16'd20;
        RAM_0[450] = -16'd3;
        RAM_1[450] = 16'd2;
        RAM_2[450] = -16'd11;
        RAM_3[450] = 16'd12;
        RAM_0[451] = -16'd2;
        RAM_1[451] = -16'd11;
        RAM_2[451] = -16'd4;
        RAM_3[451] = 16'd5;
        RAM_0[452] = -16'd6;
        RAM_1[452] = 16'd0;
        RAM_2[452] = 16'd0;
        RAM_3[452] = 16'd0;
        RAM_0[453] = -16'd1;
        RAM_1[453] = -16'd3;
        RAM_2[453] = -16'd8;
        RAM_3[453] = -16'd8;
        RAM_0[454] = 16'd1;
        RAM_1[454] = -16'd20;
        RAM_2[454] = -16'd24;
        RAM_3[454] = 16'd4;
        RAM_0[455] = -16'd3;
        RAM_1[455] = -16'd2;
        RAM_2[455] = -16'd16;
        RAM_3[455] = 16'd12;
        RAM_0[456] = -16'd10;
        RAM_1[456] = -16'd14;
        RAM_2[456] = 16'd28;
        RAM_3[456] = 16'd10;
        RAM_0[457] = 16'd8;
        RAM_1[457] = -16'd3;
        RAM_2[457] = -16'd9;
        RAM_3[457] = 16'd1;
        RAM_0[458] = -16'd9;
        RAM_1[458] = 16'd0;
        RAM_2[458] = 16'd0;
        RAM_3[458] = 16'd0;
        RAM_0[459] = 16'd1;
        RAM_1[459] = 16'd2;
        RAM_2[459] = -16'd18;
        RAM_3[459] = 16'd13;
        RAM_0[460] = -16'd16;
        RAM_1[460] = 16'd0;
        RAM_2[460] = 16'd0;
        RAM_3[460] = 16'd0;
        RAM_0[461] = -16'd19;
        RAM_1[461] = 16'd9;
        RAM_2[461] = 16'd14;
        RAM_3[461] = 16'd7;
        RAM_0[462] = -16'd10;
        RAM_1[462] = 16'd0;
        RAM_2[462] = 16'd0;
        RAM_3[462] = 16'd0;
        RAM_0[463] = -16'd4;
        RAM_1[463] = 16'd0;
        RAM_2[463] = 16'd0;
        RAM_3[463] = 16'd0;
        RAM_0[464] = -16'd29;
        RAM_1[464] = 16'd17;
        RAM_2[464] = 16'd1;
        RAM_3[464] = -16'd1;
        RAM_0[465] = 16'd5;
        RAM_1[465] = -16'd3;
        RAM_2[465] = -16'd13;
        RAM_3[465] = -16'd2;
        RAM_0[466] = -16'd1;
        RAM_1[466] = 16'd4;
        RAM_2[466] = -16'd9;
        RAM_3[466] = 16'd19;
        RAM_0[467] = 16'd0;
        RAM_1[467] = -16'd8;
        RAM_2[467] = 16'd14;
        RAM_3[467] = 16'd10;
        RAM_0[468] = 16'd1;
        RAM_1[468] = -16'd20;
        RAM_2[468] = -16'd32;
        RAM_3[468] = 16'd3;
        RAM_0[469] = 16'd7;
        RAM_1[469] = -16'd10;
        RAM_2[469] = -16'd7;
        RAM_3[469] = -16'd6;
        RAM_0[470] = 16'd4;
        RAM_1[470] = -16'd9;
        RAM_2[470] = -16'd11;
        RAM_3[470] = 16'd19;
        RAM_0[471] = -16'd5;
        RAM_1[471] = -16'd5;
        RAM_2[471] = 16'd4;
        RAM_3[471] = 16'd1;
        RAM_0[472] = 16'd1;
        RAM_1[472] = 16'd0;
        RAM_2[472] = 16'd3;
        RAM_3[472] = 16'd7;
        RAM_0[473] = 16'd8;
        RAM_1[473] = -16'd13;
        RAM_2[473] = -16'd12;
        RAM_3[473] = 16'd1;
        RAM_0[474] = 16'd6;
        RAM_1[474] = -16'd12;
        RAM_2[474] = -16'd8;
        RAM_3[474] = 16'd8;
        RAM_0[475] = 16'd0;
        RAM_1[475] = 16'd1;
        RAM_2[475] = 16'd4;
        RAM_3[475] = 16'd12;
        RAM_0[476] = 16'd2;
        RAM_1[476] = -16'd4;
        RAM_2[476] = -16'd9;
        RAM_3[476] = 16'd23;
        RAM_0[477] = -16'd3;
        RAM_1[477] = -16'd15;
        RAM_2[477] = 16'd1;
        RAM_3[477] = 16'd9;
        RAM_0[478] = -16'd20;
        RAM_1[478] = -16'd4;
        RAM_2[478] = -16'd2;
        RAM_3[478] = 16'd1;
        RAM_0[479] = -16'd11;
        RAM_1[479] = 16'd0;
        RAM_2[479] = 16'd0;
        RAM_3[479] = 16'd0;
        RAM_0[480] = -16'd6;
        RAM_1[480] = 16'd37;
        RAM_2[480] = 16'd22;
        RAM_3[480] = 16'd0;
        RAM_0[481] = -16'd1;
        RAM_1[481] = 16'd14;
        RAM_2[481] = 16'd3;
        RAM_3[481] = 16'd10;
        RAM_0[482] = -16'd3;
        RAM_1[482] = 16'd18;
        RAM_2[482] = -16'd6;
        RAM_3[482] = 16'd9;
        RAM_0[483] = -16'd2;
        RAM_1[483] = 16'd8;
        RAM_2[483] = 16'd7;
        RAM_3[483] = 16'd8;
        RAM_0[484] = -16'd6;
        RAM_1[484] = 16'd0;
        RAM_2[484] = 16'd0;
        RAM_3[484] = 16'd0;
        RAM_0[485] = -16'd1;
        RAM_1[485] = -16'd25;
        RAM_2[485] = -16'd9;
        RAM_3[485] = -16'd38;
        RAM_0[486] = 16'd1;
        RAM_1[486] = 16'd20;
        RAM_2[486] = 16'd7;
        RAM_3[486] = 16'd4;
        RAM_0[487] = -16'd3;
        RAM_1[487] = 16'd23;
        RAM_2[487] = -16'd5;
        RAM_3[487] = 16'd20;
        RAM_0[488] = -16'd10;
        RAM_1[488] = -16'd14;
        RAM_2[488] = 16'd0;
        RAM_3[488] = -16'd9;
        RAM_0[489] = 16'd8;
        RAM_1[489] = -16'd5;
        RAM_2[489] = 16'd0;
        RAM_3[489] = 16'd6;
        RAM_0[490] = -16'd9;
        RAM_1[490] = 16'd0;
        RAM_2[490] = 16'd0;
        RAM_3[490] = 16'd0;
        RAM_0[491] = 16'd1;
        RAM_1[491] = 16'd14;
        RAM_2[491] = 16'd5;
        RAM_3[491] = 16'd14;
        RAM_0[492] = -16'd16;
        RAM_1[492] = 16'd0;
        RAM_2[492] = 16'd0;
        RAM_3[492] = 16'd0;
        RAM_0[493] = -16'd19;
        RAM_1[493] = -16'd6;
        RAM_2[493] = -16'd13;
        RAM_3[493] = 16'd15;
        RAM_0[494] = -16'd10;
        RAM_1[494] = 16'd0;
        RAM_2[494] = 16'd0;
        RAM_3[494] = 16'd0;
        RAM_0[495] = -16'd4;
        RAM_1[495] = 16'd0;
        RAM_2[495] = 16'd0;
        RAM_3[495] = 16'd0;
        RAM_0[496] = -16'd29;
        RAM_1[496] = -16'd14;
        RAM_2[496] = 16'd3;
        RAM_3[496] = 16'd3;
        RAM_0[497] = 16'd5;
        RAM_1[497] = -16'd8;
        RAM_2[497] = -16'd1;
        RAM_3[497] = 16'd4;
        RAM_0[498] = -16'd1;
        RAM_1[498] = 16'd11;
        RAM_2[498] = -16'd3;
        RAM_3[498] = 16'd20;
        RAM_0[499] = 16'd0;
        RAM_1[499] = -16'd19;
        RAM_2[499] = -16'd5;
        RAM_3[499] = -16'd9;
        RAM_0[500] = 16'd1;
        RAM_1[500] = 16'd7;
        RAM_2[500] = -16'd6;
        RAM_3[500] = 16'd5;
        RAM_0[501] = 16'd7;
        RAM_1[501] = -16'd20;
        RAM_2[501] = -16'd8;
        RAM_3[501] = 16'd2;
        RAM_0[502] = 16'd4;
        RAM_1[502] = 16'd15;
        RAM_2[502] = -16'd2;
        RAM_3[502] = 16'd2;
        RAM_0[503] = -16'd5;
        RAM_1[503] = -16'd34;
        RAM_2[503] = -16'd1;
        RAM_3[503] = -16'd13;
        RAM_0[504] = 16'd1;
        RAM_1[504] = 16'd1;
        RAM_2[504] = 16'd3;
        RAM_3[504] = 16'd25;
        RAM_0[505] = 16'd8;
        RAM_1[505] = -16'd3;
        RAM_2[505] = -16'd1;
        RAM_3[505] = 16'd2;
        RAM_0[506] = 16'd6;
        RAM_1[506] = -16'd7;
        RAM_2[506] = -16'd6;
        RAM_3[506] = 16'd1;
        RAM_0[507] = 16'd0;
        RAM_1[507] = -16'd17;
        RAM_2[507] = -16'd5;
        RAM_3[507] = 16'd2;
        RAM_0[508] = 16'd2;
        RAM_1[508] = -16'd11;
        RAM_2[508] = -16'd9;
        RAM_3[508] = -16'd13;
        RAM_0[509] = -16'd3;
        RAM_1[509] = 16'd21;
        RAM_2[509] = 16'd11;
        RAM_3[509] = 16'd9;
        RAM_0[510] = -16'd20;
        RAM_1[510] = 16'd0;
        RAM_2[510] = 16'd6;
        RAM_3[510] = 16'd2;
        RAM_0[511] = -16'd11;
        RAM_1[511] = 16'd0;
        RAM_2[511] = 16'd0;
        RAM_3[511] = 16'd0;
    end
endmodule